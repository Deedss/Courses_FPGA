// nios.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module nios (
		input  wire [7:0]  blue_in_port,       //    blue.in_port
		output wire [7:0]  blue_out_port,      //        .out_port
		input  wire        clk_clk,            //     clk.clk
		input  wire [7:0]  green_in_port,      //   green.in_port
		output wire [7:0]  green_out_port,     //        .out_port
		input  wire [7:0]  red_in_port,        //     red.in_port
		output wire [7:0]  red_out_port,       //        .out_port
		inout  wire        sd_card_b_sd_cmd,   // sd_card.b_sd_cmd
		inout  wire        sd_card_b_sd_dat,   //        .b_sd_dat
		inout  wire        sd_card_b_sd_dat3,  //        .b_sd_dat3
		output wire        sd_card_o_sd_clock, //        .o_sd_clock
		input  wire [17:0] sw_in_port,         //      sw.in_port
		output wire [17:0] sw_out_port         //        .out_port
	);

	wire          altpll_0_c0_clk;                                                                        // altpll_0:c0 -> [Altera_UP_SD_Card_Avalon_Interface_0:i_clock, SW:clk, blue:clk, green:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, red:clk, rst_controller:clk]
	wire          nios2_gen2_0_debug_reset_request_reset;                                                 // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [31:0] nios2_gen2_0_data_master_readdata;                                                      // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                                                   // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                                                   // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire   [16:0] nios2_gen2_0_data_master_address;                                                       // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                                                    // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                                                          // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_write;                                                         // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                                                     // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                                               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                                            // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [16:0] nios2_gen2_0_instruction_master_address;                                                // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                                                   // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                               // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                            // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire          mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire   [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata;    // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	wire          mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest; // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	wire    [7:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address;     // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire          mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read;        // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire    [3:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire          mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write;       // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire   [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata;   // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                                // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                             // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                                          // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire    [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                           // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire          mm_interconnect_0_altpll_0_pll_slave_read;                                              // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire          mm_interconnect_0_altpll_0_pll_slave_write;                                             // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire   [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                                         // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire          mm_interconnect_0_sw_s1_chipselect;                                                     // mm_interconnect_0:SW_s1_chipselect -> SW:chipselect
	wire   [31:0] mm_interconnect_0_sw_s1_readdata;                                                       // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire    [1:0] mm_interconnect_0_sw_s1_address;                                                        // mm_interconnect_0:SW_s1_address -> SW:address
	wire          mm_interconnect_0_sw_s1_write;                                                          // mm_interconnect_0:SW_s1_write -> SW:write_n
	wire   [31:0] mm_interconnect_0_sw_s1_writedata;                                                      // mm_interconnect_0:SW_s1_writedata -> SW:writedata
	wire          mm_interconnect_0_blue_s1_chipselect;                                                   // mm_interconnect_0:blue_s1_chipselect -> blue:chipselect
	wire   [31:0] mm_interconnect_0_blue_s1_readdata;                                                     // blue:readdata -> mm_interconnect_0:blue_s1_readdata
	wire    [1:0] mm_interconnect_0_blue_s1_address;                                                      // mm_interconnect_0:blue_s1_address -> blue:address
	wire          mm_interconnect_0_blue_s1_write;                                                        // mm_interconnect_0:blue_s1_write -> blue:write_n
	wire   [31:0] mm_interconnect_0_blue_s1_writedata;                                                    // mm_interconnect_0:blue_s1_writedata -> blue:writedata
	wire          mm_interconnect_0_green_s1_chipselect;                                                  // mm_interconnect_0:green_s1_chipselect -> green:chipselect
	wire   [31:0] mm_interconnect_0_green_s1_readdata;                                                    // green:readdata -> mm_interconnect_0:green_s1_readdata
	wire    [1:0] mm_interconnect_0_green_s1_address;                                                     // mm_interconnect_0:green_s1_address -> green:address
	wire          mm_interconnect_0_green_s1_write;                                                       // mm_interconnect_0:green_s1_write -> green:write_n
	wire   [31:0] mm_interconnect_0_green_s1_writedata;                                                   // mm_interconnect_0:green_s1_writedata -> green:writedata
	wire          mm_interconnect_0_red_s1_chipselect;                                                    // mm_interconnect_0:red_s1_chipselect -> red:chipselect
	wire   [31:0] mm_interconnect_0_red_s1_readdata;                                                      // red:readdata -> mm_interconnect_0:red_s1_readdata
	wire    [1:0] mm_interconnect_0_red_s1_address;                                                       // mm_interconnect_0:red_s1_address -> red:address
	wire          mm_interconnect_0_red_s1_write;                                                         // mm_interconnect_0:red_s1_write -> red:write_n
	wire   [31:0] mm_interconnect_0_red_s1_writedata;                                                     // mm_interconnect_0:red_s1_writedata -> red:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                       // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [127:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                         // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [10:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                          // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [15:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                       // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                                            // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [127:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                        // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                                            // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          irq_mapper_receiver0_irq;                                                               // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] nios2_gen2_0_irq_irq;                                                                   // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire          rst_controller_reset_out_reset;                                                         // rst_controller:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, SW:reset_n, blue:reset_n, green:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, red:reset_n, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                                                     // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                                     // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (altpll_0_c0_clk),                                                                        //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                                        //               reset.reset_n
		.b_SD_cmd             (sd_card_b_sd_cmd),                                                                       //         conduit_end.b_sd_cmd
		.b_SD_dat             (sd_card_b_sd_dat),                                                                       //                    .b_sd_dat
		.b_SD_dat3            (sd_card_b_sd_dat3),                                                                      //                    .b_sd_dat3
		.o_SD_clock           (sd_card_o_sd_clock)                                                                      //                    .o_sd_clock
	);

	nios_SW sw (
		.clk        (altpll_0_c0_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_in_port),                         // external_connection.export
		.out_port   (sw_out_port)                         //                    .export
	);

	nios_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	nios_blue blue (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_blue_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_blue_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_blue_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_blue_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_blue_s1_readdata),   //                    .readdata
		.in_port    (blue_in_port),                         // external_connection.export
		.out_port   (blue_out_port)                         //                    .export
	);

	nios_green green (
		.clk        (altpll_0_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_s1_readdata),   //                    .readdata
		.in_port    (green_in_port),                         // external_connection.export
		.out_port   (green_out_port)                         //                    .export
	);

	nios_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_green red (
		.clk        (altpll_0_c0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_s1_readdata),   //                    .readdata
		.in_port    (red_in_port),                         // external_connection.export
		.out_port   (red_out_port)                         //                    .export
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                                      (altpll_0_c0_clk),                                                                        //                                              altpll_0_c0.clk
		.clk_0_clk_clk                                                        (clk_clk),                                                                                //                                                clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                                                     //     altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                                                         //                 nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                                     (nios2_gen2_0_data_master_address),                                                       //                                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                                 (nios2_gen2_0_data_master_waitrequest),                                                   //                                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable                                  (nios2_gen2_0_data_master_byteenable),                                                    //                                                         .byteenable
		.nios2_gen2_0_data_master_read                                        (nios2_gen2_0_data_master_read),                                                          //                                                         .read
		.nios2_gen2_0_data_master_readdata                                    (nios2_gen2_0_data_master_readdata),                                                      //                                                         .readdata
		.nios2_gen2_0_data_master_write                                       (nios2_gen2_0_data_master_write),                                                         //                                                         .write
		.nios2_gen2_0_data_master_writedata                                   (nios2_gen2_0_data_master_writedata),                                                     //                                                         .writedata
		.nios2_gen2_0_data_master_debugaccess                                 (nios2_gen2_0_data_master_debugaccess),                                                   //                                                         .debugaccess
		.nios2_gen2_0_instruction_master_address                              (nios2_gen2_0_instruction_master_address),                                                //                          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                          (nios2_gen2_0_instruction_master_waitrequest),                                            //                                                         .waitrequest
		.nios2_gen2_0_instruction_master_read                                 (nios2_gen2_0_instruction_master_read),                                                   //                                                         .read
		.nios2_gen2_0_instruction_master_readdata                             (nios2_gen2_0_instruction_master_readdata),                                               //                                                         .readdata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                                                         .write
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                                                         .read
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                                                         .readdata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                                                         .writedata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                                                         .byteenable
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                                                         .waitrequest
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  //                                                         .chipselect
		.altpll_0_pll_slave_address                                           (mm_interconnect_0_altpll_0_pll_slave_address),                                           //                                       altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                             (mm_interconnect_0_altpll_0_pll_slave_write),                                             //                                                         .write
		.altpll_0_pll_slave_read                                              (mm_interconnect_0_altpll_0_pll_slave_read),                                              //                                                         .read
		.altpll_0_pll_slave_readdata                                          (mm_interconnect_0_altpll_0_pll_slave_readdata),                                          //                                                         .readdata
		.altpll_0_pll_slave_writedata                                         (mm_interconnect_0_altpll_0_pll_slave_writedata),                                         //                                                         .writedata
		.blue_s1_address                                                      (mm_interconnect_0_blue_s1_address),                                                      //                                                  blue_s1.address
		.blue_s1_write                                                        (mm_interconnect_0_blue_s1_write),                                                        //                                                         .write
		.blue_s1_readdata                                                     (mm_interconnect_0_blue_s1_readdata),                                                     //                                                         .readdata
		.blue_s1_writedata                                                    (mm_interconnect_0_blue_s1_writedata),                                                    //                                                         .writedata
		.blue_s1_chipselect                                                   (mm_interconnect_0_blue_s1_chipselect),                                                   //                                                         .chipselect
		.green_s1_address                                                     (mm_interconnect_0_green_s1_address),                                                     //                                                 green_s1.address
		.green_s1_write                                                       (mm_interconnect_0_green_s1_write),                                                       //                                                         .write
		.green_s1_readdata                                                    (mm_interconnect_0_green_s1_readdata),                                                    //                                                         .readdata
		.green_s1_writedata                                                   (mm_interconnect_0_green_s1_writedata),                                                   //                                                         .writedata
		.green_s1_chipselect                                                  (mm_interconnect_0_green_s1_chipselect),                                                  //                                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                                //                            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                                  //                                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                   //                                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                               //                                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                              //                                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                            //                                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                             //                                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address                                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                                 //                             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                                   //                                                         .write
		.nios2_gen2_0_debug_mem_slave_read                                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                                    //                                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                                //                                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                               //                                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),                              //                                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),                             //                                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),                             //                                                         .debugaccess
		.onchip_memory2_0_s1_address                                          (mm_interconnect_0_onchip_memory2_0_s1_address),                                          //                                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                            (mm_interconnect_0_onchip_memory2_0_s1_write),                                            //                                                         .write
		.onchip_memory2_0_s1_readdata                                         (mm_interconnect_0_onchip_memory2_0_s1_readdata),                                         //                                                         .readdata
		.onchip_memory2_0_s1_writedata                                        (mm_interconnect_0_onchip_memory2_0_s1_writedata),                                        //                                                         .writedata
		.onchip_memory2_0_s1_byteenable                                       (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                                       //                                                         .byteenable
		.onchip_memory2_0_s1_chipselect                                       (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                                       //                                                         .chipselect
		.onchip_memory2_0_s1_clken                                            (mm_interconnect_0_onchip_memory2_0_s1_clken),                                            //                                                         .clken
		.red_s1_address                                                       (mm_interconnect_0_red_s1_address),                                                       //                                                   red_s1.address
		.red_s1_write                                                         (mm_interconnect_0_red_s1_write),                                                         //                                                         .write
		.red_s1_readdata                                                      (mm_interconnect_0_red_s1_readdata),                                                      //                                                         .readdata
		.red_s1_writedata                                                     (mm_interconnect_0_red_s1_writedata),                                                     //                                                         .writedata
		.red_s1_chipselect                                                    (mm_interconnect_0_red_s1_chipselect),                                                    //                                                         .chipselect
		.SW_s1_address                                                        (mm_interconnect_0_sw_s1_address),                                                        //                                                    SW_s1.address
		.SW_s1_write                                                          (mm_interconnect_0_sw_s1_write),                                                          //                                                         .write
		.SW_s1_readdata                                                       (mm_interconnect_0_sw_s1_readdata),                                                       //                                                         .readdata
		.SW_s1_writedata                                                      (mm_interconnect_0_sw_s1_writedata),                                                      //                                                         .writedata
		.SW_s1_chipselect                                                     (mm_interconnect_0_sw_s1_chipselect)                                                      //                                                         .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
