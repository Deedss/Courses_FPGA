module colourfiltering(

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK_50,

	//////////// LED //////////
	output		     [8:0]		LEDG,
	output		    [17:0]		LEDR,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,
	output		     [6:0]		HEX6,
	output		     [6:0]		HEX7,
	
	//////////// SW //////////
	input 		    [17:0]		SW,

	//////////// SD //////////
	inout   			SD_DAT, 
	inout   			SD_CMD, 
	inout   			SD_DAT3, 
	output  			SD_CLOCK,	

	//////////// RS232 //////////
	input 		          		UART_CTS,
	output		          		UART_RTS,
	input 		          		UART_RXD,
	output		          		UART_TXD,

	//////////// VGA //////////
	output		          		VGA_BLANK_N,
	output		     [7:0]		VGA_B,
	output		          		VGA_CLK,
	output		     [7:0]		VGA_G,
	output		          		VGA_HS,
	output		     [7:0]		VGA_R,
	output		          		VGA_SYNC_N,
	output		          		VGA_VS,

	//////////// GPIO, GPIO connect to D8M-GPIO //////////
	inout 		          		CAMERA_I2C_SCL,
	inout 		          		CAMERA_I2C_SDA,
	output		          		CAMERA_PWDN_n,
	output		          		MIPI_CS_n,
	inout 		          		MIPI_I2C_SCL,
	inout 		          		MIPI_I2C_SDA,
	output		          		MIPI_MCLK,
	input 		          		MIPI_PIXEL_CLK,
	input 		     [9:0]		MIPI_PIXEL_D,
	input 		          		MIPI_PIXEL_HS,
	input 		          		MIPI_PIXEL_VS,
	output		          		MIPI_REFCLK,
	output		          		MIPI_RESET_n
);

//=============================================================================
// REG/WIRE declarations
//=============================================================================
  wire        AUTO_FOC ;
  wire        READ_Request ;
  wire 	[7:0]VGA_B_A;
  wire 	[7:0]VGA_G_A;
  wire 	[7:0]VGA_R_A;
  wire        VGA_CLK_25M ;
  wire        RESET_N  ; 
  wire  [7:0]sCCD_R;
  wire  [7:0]sCCD_G;
  wire  [7:0]sCCD_B; 
  wire [15:0] H_Cont ; 
  wire [15:0] V_Cont ; 
  wire        I2C_RELEASE ;  
  wire        CAMERA_I2C_SCL_MIPI ; 
  wire        CAMERA_I2C_SCL_AF ;
  wire        CAMERA_MIPI_RELAESE ;
  wire        MIPI_BRIDGE_RELEASE ;
  wire        D8M_CK_HZ  ; 
  wire        D8M_CK_HZ2 ; 
  wire        D8M_CK_HZ3 ; 
  wire        RESET_KEY ; 
  wire   [9:0]MIPI_PIXEL_D_ ;
  wire        MIPI_PIXEL_VS_; 
  wire        MIPI_PIXEL_HS_;  
  
wire        LUT_MIPI_PIXEL_HS;
wire        LUT_MIPI_PIXEL_VS;
wire [9:0]  LUT_MIPI_PIXEL_D  ;
wire        MIPI_PIXEL_CLK_; 
//=======================================================
// Structural coding
//=======================================================

//--INPU MIPI-PIXEL-CLOCK DELAY
CLOCK_DELAY  del1(  .iCLK (MIPI_PIXEL_CLK),  .oCLK (MIPI_PIXEL_CLK_ ) );

//--D8M INPUT Gamma Correction              
 D8M_LUT  g_lut(
	.enable           (0) , // SW[0]            ),
	.PIXEL_CLK        (MIPI_PIXEL_CLK_   ),
	.MIPI_PIXEL_HS    (MIPI_PIXEL_HS    ),
	.MIPI_PIXEL_VS    (MIPI_PIXEL_VS    ),
	.MIPI_PIXEL_D     (MIPI_PIXEL_D     ),
	.NEW_MIPI_PIXEL_HS(LUT_MIPI_PIXEL_HS),
	.NEW_MIPI_PIXEL_VS(LUT_MIPI_PIXEL_VS),
	.NEW_MIPI_PIXEL_D (LUT_MIPI_PIXEL_D )
);




assign UART_RTS =0; 
assign UART_TXD =0; 
assign RESET_KEY      = KEY[0]; 

//----- RESET RELAY  --		
RESET_DELAY			u2	(	
							.iRST  ( RESET_KEY ),
                     .iCLK  ( CLOCK2_50 ),				
						   .oREADY( RESET_N)  
							
						);

assign MIPI_RESET_n   = RESET_N;
assign CAMERA_PWDN_n  = RESET_KEY; 
assign MIPI_CS_n      = 0; 

//------ CAMERA I2C COM BUS --------------------
assign I2C_RELEASE    = CAMERA_MIPI_RELAESE & MIPI_BRIDGE_RELEASE; 
assign CAMERA_I2C_SCL = ( I2C_RELEASE  )? CAMERA_I2C_SCL_AF  : CAMERA_I2C_SCL_MIPI ;   
 
//------ MIPI BRIDGE  I2C SETTING--------------- 
MIPI_BRIDGE_CAMERA_Config    cfin(
   .RESET_N           ( RESET_N  ), 
   .CLK_50            ( CLOCK2_50), 
   .MIPI_I2C_SCL      ( MIPI_I2C_SCL ), 
   .MIPI_I2C_SDA      ( MIPI_I2C_SDA ), 
   .MIPI_I2C_RELEASE  ( MIPI_BRIDGE_RELEASE ),  
   .CAMERA_I2C_SCL    ( CAMERA_I2C_SCL_MIPI ),
   .CAMERA_I2C_SDA    ( CAMERA_I2C_SDA ),
   .CAMERA_I2C_RELAESE( CAMERA_MIPI_RELAESE )
);
 
//-- Video PLL --- 
pll_test  ref(
	   .inclk0    ( CLOCK2_50 ),
	   .areset       ( 1'b0 ),
	   .c0  ( MIPI_REFCLK ),    //20Mhz
	   .c1  ( VGA_CLK_25M )    //25Mhz
		);

//--- D8M RAWDATA to RGB ---
D8M_SET   ccd (
	.RESET_SYS_N  ( RESET_N ),
   .CLOCK_50     ( CLOCK2_50      ),
	.CCD_DATA     ( LUT_MIPI_PIXEL_D [9:0]) ,
	.CCD_FVAL     ( LUT_MIPI_PIXEL_VS ), //60HZ
	.CCD_LVAL	  ( LUT_MIPI_PIXEL_HS ), // 
	.CCD_PIXCLK   ( MIPI_PIXEL_CLK_), //25MHZ
	.READ_EN      (READ_Request) , 	
   .VGA_CLK      ( VGA_CLK),
   .VGA_HS       ( VGA_HS ),
   .VGA_VS       ( VGA_VS ),	
	.X_Cont       ( H_Cont),  
   .Y_Cont       ( V_Cont),   
   .sCCD_R       ( sCCD_R ),
   .sCCD_G       ( sCCD_G ),
   .sCCD_B       ( sCCD_B )
);

//--- By Trigged VGA Controller --  
VGA_Controller_trig	u1	(
	  .iCLK       ( VGA_CLK_25M ), 
     .H_Cont		(H_Cont),  
     .V_Cont		(V_Cont),  
	  .READ_Request(READ_Request)	 , 	  
     .iRed       ( sCCD_R ),
	  .iGreen     ( sCCD_G  ),
	  .iBlue      ( sCCD_B ),		
	  .oVGA_R     ( VGA_R_A ),
	  .oVGA_G     ( VGA_G_A ),
	  .oVGA_B     ( VGA_B_A ),
     .oVGA_H_SYNC( VGA_HS ),
     .oVGA_V_SYNC( VGA_VS ),	  
	  .oVGA_SYNC  ( VGA_SYNC_N  ),
	  .oVGA_BLANK ( VGA_BLANK_N ),
	  .oVGA_CLOCK ( VGA_CLK     ),
	  .iRST_N     ( RESET_N )	
);

					
nios nios1(
	.clk_clk 			(CLOCK_50),   				// clk.clk
	.blue_in_port		(VGA_B_A), 				// blue.in_port
	.blue_out_port		(VGA_B),  				// .out_port
	.green_in_port		(VGA_G_A), 				// green.in_port
	.green_out_port	(VGA_G), 				// .out_port
	.red_in_port		(VGA_R_A), 					// red.in_port
	.red_out_port    	(VGA_R),				// .out_port
	.sw_in_port			(SW[17:0]),				// SWITCHES
	.sw_out_port		(LEDR[17:0]),			// LEDR
	.sd_card_b_sd_cmd	(SD_CMD),   // sd_card.b_sd_cmd
	.sd_card_b_sd_dat	(SD_DAT),   //        .b_sd_dat
	.sd_card_b_sd_dat3(SD_DAT3),  //        .b_sd_dat3
	.sd_card_o_sd_clock	(SD_CLK), //        .o_sd_clock
);								  
								  

//--Frame Counter -- 
 FpsMonitor uFps2(
	  .clk50    ( CLOCK2_50 ),
	  .vs       ( VGA_VS    ),//LUT_MIPI_PIXEL_VS ), //60HZ
	  .fps      (  ),
	  .hex_fps_h( HEX1 ),
	  .hex_fps_l( HEX0 )
);

////----7-SEG OFF----
assign  HEX2 = 7'h7F;
assign  HEX3 = 7'h7F;
assign  HEX4 = 7'h7F;
assign  HEX5 = 7'h7F;
assign  HEX6 = 7'h7F;
assign  HEX7 = 7'h7F;

//--FREQUNCY TEST--
CLOCKMEM  ck1 ( .CLK(VGA_CLK_25M    ),.CLK_FREQ  (25000000  ),.CK_1HZ (D8M_CK_HZ   ));
CLOCKMEM  ck2 ( .CLK(MIPI_REFCLK    ),.CLK_FREQ  (20000000  ),.CK_1HZ (D8M_CK_HZ2  ));
CLOCKMEM  ck3 ( .CLK(MIPI_PIXEL_CLK_),.CLK_FREQ  (25000000 ),.CK_1HZ (D8M_CK_HZ3   ));

//--LED STATUS-----
//assign LEDR[9:0] = { D8M_CK_HZ ,D8M_CK_HZ2,D8M_CK_HZ3 ,5'h0,CAMERA_MIPI_RELAESE ,MIPI_BRIDGE_RELEASE } ; 
endmodule
