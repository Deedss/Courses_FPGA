// nios.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module nios (
		input  wire        clk_clk,       //     clk.clk
		input  wire        reset_reset_n, //   reset.reset_n
		inout  wire [15:0] sram_DQ,       //    sram.DQ
		output wire [19:0] sram_ADDR,     //        .ADDR
		output wire        sram_LB_N,     //        .LB_N
		output wire        sram_UB_N,     //        .UB_N
		output wire        sram_CE_N,     //        .CE_N
		output wire        sram_OE_N,     //        .OE_N
		output wire        sram_WE_N,     //        .WE_N
		output wire        vga_out_CLK,   // vga_out.CLK
		output wire        vga_out_HS,    //        .HS
		output wire        vga_out_VS,    //        .VS
		output wire        vga_out_BLANK, //        .BLANK
		output wire        vga_out_SYNC,  //        .SYNC
		output wire [7:0]  vga_out_R,     //        .R
		output wire [7:0]  vga_out_G,     //        .G
		output wire [7:0]  vga_out_B      //        .B
	);

	wire         video_dma_controller_0_avalon_pixel_source_valid;                             // video_dma_controller_0:stream_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dma_controller_0_avalon_pixel_source_data;                              // video_dma_controller_0:stream_data -> video_vga_controller_0:data
	wire         video_dma_controller_0_avalon_pixel_source_ready;                             // video_vga_controller_0:ready -> video_dma_controller_0:stream_ready
	wire         video_dma_controller_0_avalon_pixel_source_startofpacket;                     // video_dma_controller_0:stream_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dma_controller_0_avalon_pixel_source_endofpacket;                       // video_dma_controller_0:stream_endofpacket -> video_vga_controller_0:endofpacket
	wire         altpll_0_c0_clk;                                                              // altpll_0:c0 -> [mm_interconnect_0:altpll_0_c0_clk, rst_controller_001:clk, video_dma_controller_0:clk, video_vga_controller_0:clk]
	wire         video_dma_controller_0_avalon_dma_master_waitrequest;                         // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	wire  [31:0] video_dma_controller_0_avalon_dma_master_readdata;                            // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	wire  [31:0] video_dma_controller_0_avalon_dma_master_address;                             // video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	wire         video_dma_controller_0_avalon_dma_master_read;                                // video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	wire         video_dma_controller_0_avalon_dma_master_readdatavalid;                       // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	wire         video_dma_controller_0_avalon_dma_master_lock;                                // video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                            // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                         // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                         // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [21:0] nios2_gen2_0_data_master_address;                                             // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                          // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                                       // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                               // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                           // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                     // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                  // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [21:0] nios2_gen2_0_instruction_master_address;                                      // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                         // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                                // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_readdata;                          // sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_0_avalon_sram_slave_address;                           // mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_read;                              // mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	wire   [1:0] mm_interconnect_0_sram_0_avalon_sram_slave_byteenable;                        // mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid;                     // sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_write;                             // mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_writedata;                         // mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	wire  [31:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata;   // video_dma_controller_0:slave_readdata -> mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address;    // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	wire         mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read;       // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	wire   [3:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable; // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	wire         mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write;      // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	wire  [31:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata;  // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                      // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                   // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                                // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                 // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                                    // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                                   // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                               // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                         // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [altpll_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sram_0:reset]
	wire         rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, video_dma_controller_0:reset, video_vga_controller_0:reset]

	nios_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	nios_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_sram_0 sram_0 (
		.clk           (clk_clk),                                                  //                clk.clk
		.reset         (rst_controller_reset_out_reset),                           //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                  // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                //                   .export
		.address       (mm_interconnect_0_sram_0_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_0_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_0_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.master_address       (video_dma_controller_0_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma_controller_0_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma_controller_0_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma_controller_0_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma_controller_0_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma_controller_0_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma_controller_0_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma_controller_0_avalon_pixel_source_valid)                              //                         .valid
	);

	nios_video_vga_controller_0 video_vga_controller_0 (
		.clk           (altpll_0_c0_clk),                                          //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                       //              reset.reset
		.data          (video_dma_controller_0_avalon_pixel_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),   //                   .endofpacket
		.valid         (video_dma_controller_0_avalon_pixel_source_valid),         //                   .valid
		.ready         (video_dma_controller_0_avalon_pixel_source_ready),         //                   .ready
		.VGA_CLK       (vga_out_CLK),                                              // external_interface.export
		.VGA_HS        (vga_out_HS),                                               //                   .export
		.VGA_VS        (vga_out_VS),                                               //                   .export
		.VGA_BLANK     (vga_out_BLANK),                                            //                   .export
		.VGA_SYNC      (vga_out_SYNC),                                             //                   .export
		.VGA_R         (vga_out_R),                                                //                   .export
		.VGA_G         (vga_out_G),                                                //                   .export
		.VGA_B         (vga_out_B)                                                 //                   .export
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                                              //                                          altpll_0_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                                      //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                               // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                                           //   video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                                             //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                                         //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                                          //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                                //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                                            //                                                     .readdata
		.nios2_gen2_0_data_master_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                                       //                                                     .readdatavalid
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                               //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                                           //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                                         //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                                      //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                                  //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                                         //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                                     //                                                     .readdata
		.nios2_gen2_0_instruction_master_readdatavalid              (nios2_gen2_0_instruction_master_readdatavalid),                                //                                                     .readdatavalid
		.video_dma_controller_0_avalon_dma_master_address           (video_dma_controller_0_avalon_dma_master_address),                             //             video_dma_controller_0_avalon_dma_master.address
		.video_dma_controller_0_avalon_dma_master_waitrequest       (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                                                     .waitrequest
		.video_dma_controller_0_avalon_dma_master_read              (video_dma_controller_0_avalon_dma_master_read),                                //                                                     .read
		.video_dma_controller_0_avalon_dma_master_readdata          (video_dma_controller_0_avalon_dma_master_readdata),                            //                                                     .readdata
		.video_dma_controller_0_avalon_dma_master_readdatavalid     (video_dma_controller_0_avalon_dma_master_readdatavalid),                       //                                                     .readdatavalid
		.video_dma_controller_0_avalon_dma_master_lock              (video_dma_controller_0_avalon_dma_master_lock),                                //                                                     .lock
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                                 //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                                   //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                                    //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                                //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                               //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                      //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                        //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                         //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                     //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                    //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                  //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                   //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                       //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                         //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                          //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                      //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                     //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),                    //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),                   //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),                   //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                                //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                                  //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                               //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                              //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                             //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                             //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                                  //                                                     .clken
		.sram_0_avalon_sram_slave_address                           (mm_interconnect_0_sram_0_avalon_sram_slave_address),                           //                             sram_0_avalon_sram_slave.address
		.sram_0_avalon_sram_slave_write                             (mm_interconnect_0_sram_0_avalon_sram_slave_write),                             //                                                     .write
		.sram_0_avalon_sram_slave_read                              (mm_interconnect_0_sram_0_avalon_sram_slave_read),                              //                                                     .read
		.sram_0_avalon_sram_slave_readdata                          (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),                          //                                                     .readdata
		.sram_0_avalon_sram_slave_writedata                         (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),                         //                                                     .writedata
		.sram_0_avalon_sram_slave_byteenable                        (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),                        //                                                     .byteenable
		.sram_0_avalon_sram_slave_readdatavalid                     (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid),                     //                                                     .readdatavalid
		.video_dma_controller_0_avalon_dma_control_slave_address    (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address),    //      video_dma_controller_0_avalon_dma_control_slave.address
		.video_dma_controller_0_avalon_dma_control_slave_write      (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write),      //                                                     .write
		.video_dma_controller_0_avalon_dma_control_slave_read       (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read),       //                                                     .read
		.video_dma_controller_0_avalon_dma_control_slave_readdata   (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                                                     .readdata
		.video_dma_controller_0_avalon_dma_control_slave_writedata  (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                                                     .writedata
		.video_dma_controller_0_avalon_dma_control_slave_byteenable (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable)  //                                                     .byteenable
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
