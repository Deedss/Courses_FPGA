library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity camera_in is
	port(
		
	)